`define module_name AHB2AXI_Bridge
